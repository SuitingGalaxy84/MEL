module Twiddle512 #(
    parameter TW_FF = 1
)(
    input                 clock,
    input  [8:0]          addr,
    output [15:0]         tw_re,
    output [15:0]         tw_im
);

    wire[15:0] wn_re [0:511];
    wire[15:0] wn_im [0:511];
    wire[15:0] mx_re;
    wire[15:0] mx_im;
    reg [15:0] ff_re;
    reg [15:0] ff_im;

    assign mx_re = wn_re[addr];
    assign mx_im = wn_im[addr];

    always @(posedge clock) begin
        ff_re <= mx_re;
        ff_im <= mx_im;
    end

    assign tw_re = (TW_FF) ? ff_re :  mx_re;
    assign tw_im = (TW_FF) ? ff_im :  mx_im;

    //      wn_re = cos(-2pi*n/512)          wn_im = sin(-2pi*n/512)
    assign  wn_re[ 0] = 16'h0000;   assign  wn_im[ 0] = 16'h0000;   //  0   1.000  -0.000
    assign  wn_re[ 1] = 16'h7FFE;   assign  wn_im[ 1] = 16'hFE6E;   //  1   1.000  -0.012
    assign  wn_re[ 2] = 16'h7FF6;   assign  wn_im[ 2] = 16'hFCDC;   //  2   1.000  -0.025
    assign  wn_re[ 3] = 16'h7FEA;   assign  wn_im[ 3] = 16'hFB4A;   //  3   0.999  -0.037
    assign  wn_re[ 4] = 16'h7FD9;   assign  wn_im[ 4] = 16'hF9B8;   //  4   0.999  -0.049
    assign  wn_re[ 5] = 16'h7FC2;   assign  wn_im[ 5] = 16'hF827;   //  5   0.998  -0.061
    assign  wn_re[ 6] = 16'h7FA7;   assign  wn_im[ 6] = 16'hF695;   //  6   0.997  -0.074
    assign  wn_re[ 7] = 16'h7F87;   assign  wn_im[ 7] = 16'hF505;   //  7   0.996  -0.086
    assign  wn_re[ 8] = 16'h7F62;   assign  wn_im[ 8] = 16'hF374;   //  8   0.995  -0.098
    assign  wn_re[ 9] = 16'h7F38;   assign  wn_im[ 9] = 16'hF1E4;   //  9   0.994  -0.110
    assign  wn_re[10] = 16'h7F0A;   assign  wn_im[10] = 16'hF055;   // 10   0.992  -0.122
    assign  wn_re[11] = 16'h7ED6;   assign  wn_im[11] = 16'hEEC6;   // 11   0.991  -0.135
    assign  wn_re[12] = 16'h7E9D;   assign  wn_im[12] = 16'hED38;   // 12   0.989  -0.147
    assign  wn_re[13] = 16'h7E60;   assign  wn_im[13] = 16'hEBAB;   // 13   0.987  -0.159
    assign  wn_re[14] = 16'h7E1E;   assign  wn_im[14] = 16'hEA1E;   // 14   0.985  -0.171
    assign  wn_re[15] = 16'h7DD6;   assign  wn_im[15] = 16'hE892;   // 15   0.983  -0.183
    assign  wn_re[16] = 16'h7D8A;   assign  wn_im[16] = 16'hE707;   // 16   0.981  -0.195
    assign  wn_re[17] = 16'h7D3A;   assign  wn_im[17] = 16'hE57D;   // 17   0.978  -0.207
    assign  wn_re[18] = 16'h7CE4;   assign  wn_im[18] = 16'hE3F4;   // 18   0.976  -0.219
    assign  wn_re[19] = 16'h7C89;   assign  wn_im[19] = 16'hE26D;   // 19   0.973  -0.231
    assign  wn_re[20] = 16'h7C2A;   assign  wn_im[20] = 16'hE0E6;   // 20   0.970  -0.243
    assign  wn_re[21] = 16'h7BC6;   assign  wn_im[21] = 16'hDF61;   // 21   0.967  -0.255
    assign  wn_re[22] = 16'h7B5D;   assign  wn_im[22] = 16'hDDDC;   // 22   0.964  -0.267
    assign  wn_re[23] = 16'h7AEF;   assign  wn_im[23] = 16'hDC59;   // 23   0.960  -0.279
    assign  wn_re[24] = 16'h7A7D;   assign  wn_im[24] = 16'hDAD8;   // 24   0.957  -0.290
    assign  wn_re[25] = 16'h7A06;   assign  wn_im[25] = 16'hD958;   // 25   0.953  -0.302
    assign  wn_re[26] = 16'h798A;   assign  wn_im[26] = 16'hD7D9;   // 26   0.950  -0.314
    assign  wn_re[27] = 16'h790A;   assign  wn_im[27] = 16'hD65C;   // 27   0.946  -0.325
    assign  wn_re[28] = 16'h7885;   assign  wn_im[28] = 16'hD4E1;   // 28   0.942  -0.337
    assign  wn_re[29] = 16'h77FB;   assign  wn_im[29] = 16'hD367;   // 29   0.937  -0.348
    assign  wn_re[30] = 16'h776C;   assign  wn_im[30] = 16'hD1EF;   // 30   0.933  -0.360
    assign  wn_re[31] = 16'h76D9;   assign  wn_im[31] = 16'hD079;   // 31   0.929  -0.371
    assign  wn_re[32] = 16'h7642;   assign  wn_im[32] = 16'hCF04;   // 32   0.924  -0.383
    assign  wn_re[33] = 16'h75A6;   assign  wn_im[33] = 16'hCD92;   // 33   0.919  -0.394
    assign  wn_re[34] = 16'h7505;   assign  wn_im[34] = 16'hCC21;   // 34   0.914  -0.405
    assign  wn_re[35] = 16'h7460;   assign  wn_im[35] = 16'hCAB2;   // 35   0.909  -0.416
    assign  wn_re[36] = 16'h73B6;   assign  wn_im[36] = 16'hC946;   // 36   0.904  -0.428
    assign  wn_re[37] = 16'h7308;   assign  wn_im[37] = 16'hC7DB;   // 37   0.899  -0.439
    assign  wn_re[38] = 16'h7255;   assign  wn_im[38] = 16'hC673;   // 38   0.893  -0.450
    assign  wn_re[39] = 16'h719E;   assign  wn_im[39] = 16'hC50D;   // 39   0.888  -0.461
    assign  wn_re[40] = 16'h70E3;   assign  wn_im[40] = 16'hC3A9;   // 40   0.882  -0.471
    assign  wn_re[41] = 16'h7023;   assign  wn_im[41] = 16'hC248;   // 41   0.876  -0.482
    assign  wn_re[42] = 16'h6F5F;   assign  wn_im[42] = 16'hC0E9;   // 42   0.870  -0.493
    assign  wn_re[43] = 16'h6E97;   assign  wn_im[43] = 16'hBF8C;   // 43   0.864  -0.504
    assign  wn_re[44] = 16'h6DCA;   assign  wn_im[44] = 16'hBE32;   // 44   0.858  -0.514
    assign  wn_re[45] = 16'h6CF9;   assign  wn_im[45] = 16'hBCDA;   // 45   0.851  -0.525
    assign  wn_re[46] = 16'h6C24;   assign  wn_im[46] = 16'hBB85;   // 46   0.845  -0.535
    assign  wn_re[47] = 16'h6B4B;   assign  wn_im[47] = 16'hBA33;   // 47   0.838  -0.545
    assign  wn_re[48] = 16'h6A6E;   assign  wn_im[48] = 16'hB8E3;   // 48   0.831  -0.556
    assign  wn_re[49] = 16'h698C;   assign  wn_im[49] = 16'hB796;   // 49   0.825  -0.566
    assign  wn_re[50] = 16'h68A7;   assign  wn_im[50] = 16'hB64C;   // 50   0.818  -0.576
    assign  wn_re[51] = 16'h67BD;   assign  wn_im[51] = 16'hB505;   // 51   0.810  -0.586
    assign  wn_re[52] = 16'h66D0;   assign  wn_im[52] = 16'hB3C0;   // 52   0.803  -0.596
    assign  wn_re[53] = 16'h65DE;   assign  wn_im[53] = 16'hB27F;   // 53   0.796  -0.606
    assign  wn_re[54] = 16'h64E9;   assign  wn_im[54] = 16'hB140;   // 54   0.788  -0.615
    assign  wn_re[55] = 16'h63EF;   assign  wn_im[55] = 16'hB005;   // 55   0.781  -0.625
    assign  wn_re[56] = 16'h62F2;   assign  wn_im[56] = 16'hAECC;   // 56   0.773  -0.634
    assign  wn_re[57] = 16'h61F1;   assign  wn_im[57] = 16'hAD97;   // 57   0.765  -0.644
    assign  wn_re[58] = 16'h60EC;   assign  wn_im[58] = 16'hAC65;   // 58   0.757  -0.653
    assign  wn_re[59] = 16'h5FE4;   assign  wn_im[59] = 16'hAB36;   // 59   0.749  -0.662
    assign  wn_re[60] = 16'h5ED7;   assign  wn_im[60] = 16'hAA0A;   // 60   0.741  -0.672
    assign  wn_re[61] = 16'h5DC8;   assign  wn_im[61] = 16'hA8E2;   // 61   0.733  -0.681
    assign  wn_re[62] = 16'h5CB4;   assign  wn_im[62] = 16'hA7BD;   // 62   0.724  -0.690
    assign  wn_re[63] = 16'h5B9D;   assign  wn_im[63] = 16'hA69C;   // 63   0.716  -0.698
    assign  wn_re[64] = 16'h5A82;   assign  wn_im[64] = 16'hA57E;   // 64   0.707  -0.707
    assign  wn_re[65] = 16'h5964;   assign  wn_im[65] = 16'hA463;   // 65   0.698  -0.716
    assign  wn_re[66] = 16'h5843;   assign  wn_im[66] = 16'hA34C;   // 66   0.690  -0.724
    assign  wn_re[67] = 16'h571E;   assign  wn_im[67] = 16'hA238;   // 67   0.681  -0.733
    assign  wn_re[68] = 16'h55F6;   assign  wn_im[68] = 16'hA129;   // 68   0.672  -0.741
    assign  wn_re[69] = 16'h54CA;   assign  wn_im[69] = 16'hA01C;   // 69   0.662  -0.749
    assign  wn_re[70] = 16'h539B;   assign  wn_im[70] = 16'h9F14;   // 70   0.653  -0.757
    assign  wn_re[71] = 16'h5269;   assign  wn_im[71] = 16'h9E0F;   // 71   0.644  -0.765
    assign  wn_re[72] = 16'h5134;   assign  wn_im[72] = 16'h9D0E;   // 72   0.634  -0.773
    assign  wn_re[73] = 16'h4FFB;   assign  wn_im[73] = 16'h9C11;   // 73   0.625  -0.781
    assign  wn_re[74] = 16'h4EC0;   assign  wn_im[74] = 16'h9B17;   // 74   0.615  -0.788
    assign  wn_re[75] = 16'h4D81;   assign  wn_im[75] = 16'h9A22;   // 75   0.606  -0.796
    assign  wn_re[76] = 16'h4C40;   assign  wn_im[76] = 16'h9930;   // 76   0.596  -0.803
    assign  wn_re[77] = 16'h4AFB;   assign  wn_im[77] = 16'h9843;   // 77   0.586  -0.810
    assign  wn_re[78] = 16'h49B4;   assign  wn_im[78] = 16'h9759;   // 78   0.576  -0.818
    assign  wn_re[79] = 16'h486A;   assign  wn_im[79] = 16'h9674;   // 79   0.566  -0.825
    assign  wn_re[80] = 16'h471D;   assign  wn_im[80] = 16'h9592;   // 80   0.556  -0.831
    assign  wn_re[81] = 16'h45CD;   assign  wn_im[81] = 16'h94B5;   // 81   0.545  -0.838
    assign  wn_re[82] = 16'h447B;   assign  wn_im[82] = 16'h93DC;   // 82   0.535  -0.845
    assign  wn_re[83] = 16'h4326;   assign  wn_im[83] = 16'h9307;   // 83   0.525  -0.851
    assign  wn_re[84] = 16'h41CE;   assign  wn_im[84] = 16'h9236;   // 84   0.514  -0.858
    assign  wn_re[85] = 16'h4074;   assign  wn_im[85] = 16'h9169;   // 85   0.504  -0.864
    assign  wn_re[86] = 16'h3F17;   assign  wn_im[86] = 16'h90A1;   // 86   0.493  -0.870
    assign  wn_re[87] = 16'h3DB8;   assign  wn_im[87] = 16'h8FDD;   // 87   0.482  -0.876
    assign  wn_re[88] = 16'h3C57;   assign  wn_im[88] = 16'h8F1D;   // 88   0.471  -0.882
    assign  wn_re[89] = 16'h3AF3;   assign  wn_im[89] = 16'h8E62;   // 89   0.461  -0.888
    assign  wn_re[90] = 16'h398D;   assign  wn_im[90] = 16'h8DAB;   // 90   0.450  -0.893
    assign  wn_re[91] = 16'h3825;   assign  wn_im[91] = 16'h8CF8;   // 91   0.439  -0.899
    assign  wn_re[92] = 16'h36BA;   assign  wn_im[92] = 16'h8C4A;   // 92   0.428  -0.904
    assign  wn_re[93] = 16'h354E;   assign  wn_im[93] = 16'h8BA0;   // 93   0.416  -0.909
    assign  wn_re[94] = 16'h33DF;   assign  wn_im[94] = 16'h8AFB;   // 94   0.405  -0.914
    assign  wn_re[95] = 16'h326E;   assign  wn_im[95] = 16'h8A5A;   // 95   0.394  -0.919
    assign  wn_re[96] = 16'h30FC;   assign  wn_im[96] = 16'h89BE;   // 96   0.383  -0.924
    assign  wn_re[97] = 16'h2F87;   assign  wn_im[97] = 16'h8927;   // 97   0.371  -0.929
    assign  wn_re[98] = 16'h2E11;   assign  wn_im[98] = 16'h8894;   // 98   0.360  -0.933
    assign  wn_re[99] = 16'h2C99;   assign  wn_im[99] = 16'h8805;   // 99   0.348  -0.937
    assign  wn_re[100] = 16'h2B1F;   assign  wn_im[100] = 16'h877B;   // 100   0.337  -0.942
    assign  wn_re[101] = 16'h29A4;   assign  wn_im[101] = 16'h86F6;   // 101   0.325  -0.946
    assign  wn_re[102] = 16'h2827;   assign  wn_im[102] = 16'h8676;   // 102   0.314  -0.950
    assign  wn_re[103] = 16'h26A8;   assign  wn_im[103] = 16'h85FA;   // 103   0.302  -0.953
    assign  wn_re[104] = 16'h2528;   assign  wn_im[104] = 16'h8583;   // 104   0.290  -0.957
    assign  wn_re[105] = 16'h23A7;   assign  wn_im[105] = 16'h8511;   // 105   0.279  -0.960
    assign  wn_re[106] = 16'h2224;   assign  wn_im[106] = 16'h84A3;   // 106   0.267  -0.964
    assign  wn_re[107] = 16'h209F;   assign  wn_im[107] = 16'h843A;   // 107   0.255  -0.967
    assign  wn_re[108] = 16'h1F1A;   assign  wn_im[108] = 16'h83D6;   // 108   0.243  -0.970
    assign  wn_re[109] = 16'h1D93;   assign  wn_im[109] = 16'h8377;   // 109   0.231  -0.973
    assign  wn_re[110] = 16'h1C0C;   assign  wn_im[110] = 16'h831C;   // 110   0.219  -0.976
    assign  wn_re[111] = 16'h1A83;   assign  wn_im[111] = 16'h82C6;   // 111   0.207  -0.978
    assign  wn_re[112] = 16'h18F9;   assign  wn_im[112] = 16'h8276;   // 112   0.195  -0.981
    assign  wn_re[113] = 16'h176E;   assign  wn_im[113] = 16'h822A;   // 113   0.183  -0.983
    assign  wn_re[114] = 16'h15E2;   assign  wn_im[114] = 16'h81E2;   // 114   0.171  -0.985
    assign  wn_re[115] = 16'h1455;   assign  wn_im[115] = 16'h81A0;   // 115   0.159  -0.987
    assign  wn_re[116] = 16'h12C8;   assign  wn_im[116] = 16'h8163;   // 116   0.147  -0.989
    assign  wn_re[117] = 16'h113A;   assign  wn_im[117] = 16'h812A;   // 117   0.135  -0.991
    assign  wn_re[118] = 16'h0FAB;   assign  wn_im[118] = 16'h80F6;   // 118   0.122  -0.992
    assign  wn_re[119] = 16'h0E1C;   assign  wn_im[119] = 16'h80C8;   // 119   0.110  -0.994
    assign  wn_re[120] = 16'h0C8C;   assign  wn_im[120] = 16'h809E;   // 120   0.098  -0.995
    assign  wn_re[121] = 16'h0AFB;   assign  wn_im[121] = 16'h8079;   // 121   0.086  -0.996
    assign  wn_re[122] = 16'h096B;   assign  wn_im[122] = 16'h8059;   // 122   0.074  -0.997
    assign  wn_re[123] = 16'h07D9;   assign  wn_im[123] = 16'h803E;   // 123   0.061  -0.998
    assign  wn_re[124] = 16'h0648;   assign  wn_im[124] = 16'h8027;   // 124   0.049  -0.999
    assign  wn_re[125] = 16'h04B6;   assign  wn_im[125] = 16'h8016;   // 125   0.037  -0.999
    assign  wn_re[126] = 16'h0324;   assign  wn_im[126] = 16'h800A;   // 126   0.025  -1.000
    assign  wn_re[127] = 16'h0192;   assign  wn_im[127] = 16'h8002;   // 127   0.012  -1.000
    assign  wn_re[128] = 16'h0000;   assign  wn_im[128] = 16'h8000;   // 128   0.000  -1.000
    assign  wn_re[129] = 16'hFE6E;   assign  wn_im[129] = 16'h8002;   // 129  -0.012  -1.000
    assign  wn_re[130] = 16'hFCDC;   assign  wn_im[130] = 16'h800A;   // 130  -0.025  -1.000
    assign  wn_re[131] = 16'hxxxx;   assign  wn_im[131] = 16'hxxxx;   // 131  -0.037  -0.999
    assign  wn_re[132] = 16'hF9B8;   assign  wn_im[132] = 16'h8027;   // 132  -0.049  -0.999
    assign  wn_re[133] = 16'hxxxx;   assign  wn_im[133] = 16'hxxxx;   // 133  -0.061  -0.998
    assign  wn_re[134] = 16'hF695;   assign  wn_im[134] = 16'h8059;   // 134  -0.074  -0.997
    assign  wn_re[135] = 16'hF505;   assign  wn_im[135] = 16'h8079;   // 135  -0.086  -0.996
    assign  wn_re[136] = 16'hF374;   assign  wn_im[136] = 16'h809E;   // 136  -0.098  -0.995
    assign  wn_re[137] = 16'hxxxx;   assign  wn_im[137] = 16'hxxxx;   // 137  -0.110  -0.994
    assign  wn_re[138] = 16'hF055;   assign  wn_im[138] = 16'h80F6;   // 138  -0.122  -0.992
    assign  wn_re[139] = 16'hxxxx;   assign  wn_im[139] = 16'hxxxx;   // 139  -0.135  -0.991
    assign  wn_re[140] = 16'hED38;   assign  wn_im[140] = 16'h8163;   // 140  -0.147  -0.989
    assign  wn_re[141] = 16'hEBAB;   assign  wn_im[141] = 16'h81A0;   // 141  -0.159  -0.987
    assign  wn_re[142] = 16'hEA1E;   assign  wn_im[142] = 16'h81E2;   // 142  -0.171  -0.985
    assign  wn_re[143] = 16'hxxxx;   assign  wn_im[143] = 16'hxxxx;   // 143  -0.183  -0.983
    assign  wn_re[144] = 16'hE707;   assign  wn_im[144] = 16'h8276;   // 144  -0.195  -0.981
    assign  wn_re[145] = 16'hxxxx;   assign  wn_im[145] = 16'hxxxx;   // 145  -0.207  -0.978
    assign  wn_re[146] = 16'hE3F4;   assign  wn_im[146] = 16'h831C;   // 146  -0.219  -0.976
    assign  wn_re[147] = 16'hE26D;   assign  wn_im[147] = 16'h8377;   // 147  -0.231  -0.973
    assign  wn_re[148] = 16'hE0E6;   assign  wn_im[148] = 16'h83D6;   // 148  -0.243  -0.970
    assign  wn_re[149] = 16'hxxxx;   assign  wn_im[149] = 16'hxxxx;   // 149  -0.255  -0.967
    assign  wn_re[150] = 16'hDDDC;   assign  wn_im[150] = 16'h84A3;   // 150  -0.267  -0.964
    assign  wn_re[151] = 16'hxxxx;   assign  wn_im[151] = 16'hxxxx;   // 151  -0.279  -0.960
    assign  wn_re[152] = 16'hDAD8;   assign  wn_im[152] = 16'h8583;   // 152  -0.290  -0.957
    assign  wn_re[153] = 16'hD958;   assign  wn_im[153] = 16'h85FA;   // 153  -0.302  -0.953
    assign  wn_re[154] = 16'hD7D9;   assign  wn_im[154] = 16'h8676;   // 154  -0.314  -0.950
    assign  wn_re[155] = 16'hxxxx;   assign  wn_im[155] = 16'hxxxx;   // 155  -0.325  -0.946
    assign  wn_re[156] = 16'hD4E1;   assign  wn_im[156] = 16'h877B;   // 156  -0.337  -0.942
    assign  wn_re[157] = 16'hxxxx;   assign  wn_im[157] = 16'hxxxx;   // 157  -0.348  -0.937
    assign  wn_re[158] = 16'hD1EF;   assign  wn_im[158] = 16'h8894;   // 158  -0.360  -0.933
    assign  wn_re[159] = 16'hD079;   assign  wn_im[159] = 16'h8927;   // 159  -0.371  -0.929
    assign  wn_re[160] = 16'hCF04;   assign  wn_im[160] = 16'h89BE;   // 160  -0.383  -0.924
    assign  wn_re[161] = 16'hxxxx;   assign  wn_im[161] = 16'hxxxx;   // 161  -0.394  -0.919
    assign  wn_re[162] = 16'hCC21;   assign  wn_im[162] = 16'h8AFB;   // 162  -0.405  -0.914
    assign  wn_re[163] = 16'hxxxx;   assign  wn_im[163] = 16'hxxxx;   // 163  -0.416  -0.909
    assign  wn_re[164] = 16'hC946;   assign  wn_im[164] = 16'h8C4A;   // 164  -0.428  -0.904
    assign  wn_re[165] = 16'hC7DB;   assign  wn_im[165] = 16'h8CF8;   // 165  -0.439  -0.899
    assign  wn_re[166] = 16'hC673;   assign  wn_im[166] = 16'h8DAB;   // 166  -0.450  -0.893
    assign  wn_re[167] = 16'hxxxx;   assign  wn_im[167] = 16'hxxxx;   // 167  -0.461  -0.888
    assign  wn_re[168] = 16'hC3A9;   assign  wn_im[168] = 16'h8F1D;   // 168  -0.471  -0.882
    assign  wn_re[169] = 16'hxxxx;   assign  wn_im[169] = 16'hxxxx;   // 169  -0.482  -0.876
    assign  wn_re[170] = 16'hC0E9;   assign  wn_im[170] = 16'h90A1;   // 170  -0.493  -0.870
    assign  wn_re[171] = 16'hBF8C;   assign  wn_im[171] = 16'h9169;   // 171  -0.504  -0.864
    assign  wn_re[172] = 16'hBE32;   assign  wn_im[172] = 16'h9236;   // 172  -0.514  -0.858
    assign  wn_re[173] = 16'hxxxx;   assign  wn_im[173] = 16'hxxxx;   // 173  -0.525  -0.851
    assign  wn_re[174] = 16'hBB85;   assign  wn_im[174] = 16'h93DC;   // 174  -0.535  -0.845
    assign  wn_re[175] = 16'hxxxx;   assign  wn_im[175] = 16'hxxxx;   // 175  -0.545  -0.838
    assign  wn_re[176] = 16'hB8E3;   assign  wn_im[176] = 16'h9592;   // 176  -0.556  -0.831
    assign  wn_re[177] = 16'hB796;   assign  wn_im[177] = 16'h9674;   // 177  -0.566  -0.825
    assign  wn_re[178] = 16'hB64C;   assign  wn_im[178] = 16'h9759;   // 178  -0.576  -0.818
    assign  wn_re[179] = 16'hxxxx;   assign  wn_im[179] = 16'hxxxx;   // 179  -0.586  -0.810
    assign  wn_re[180] = 16'hB3C0;   assign  wn_im[180] = 16'h9930;   // 180  -0.596  -0.803
    assign  wn_re[181] = 16'hxxxx;   assign  wn_im[181] = 16'hxxxx;   // 181  -0.606  -0.796
    assign  wn_re[182] = 16'hB140;   assign  wn_im[182] = 16'h9B17;   // 182  -0.615  -0.788
    assign  wn_re[183] = 16'hB005;   assign  wn_im[183] = 16'h9C11;   // 183  -0.625  -0.781
    assign  wn_re[184] = 16'hAECC;   assign  wn_im[184] = 16'h9D0E;   // 184  -0.634  -0.773
    assign  wn_re[185] = 16'hxxxx;   assign  wn_im[185] = 16'hxxxx;   // 185  -0.644  -0.765
    assign  wn_re[186] = 16'hAC65;   assign  wn_im[186] = 16'h9F14;   // 186  -0.653  -0.757
    assign  wn_re[187] = 16'hxxxx;   assign  wn_im[187] = 16'hxxxx;   // 187  -0.662  -0.749
    assign  wn_re[188] = 16'hAA0A;   assign  wn_im[188] = 16'hA129;   // 188  -0.672  -0.741
    assign  wn_re[189] = 16'hA8E2;   assign  wn_im[189] = 16'hA238;   // 189  -0.681  -0.733
    assign  wn_re[190] = 16'hA7BD;   assign  wn_im[190] = 16'hA34C;   // 190  -0.690  -0.724
    assign  wn_re[191] = 16'hxxxx;   assign  wn_im[191] = 16'hxxxx;   // 191  -0.698  -0.716
    assign  wn_re[192] = 16'hA57E;   assign  wn_im[192] = 16'hA57E;   // 192  -0.707  -0.707
    assign  wn_re[193] = 16'hxxxx;   assign  wn_im[193] = 16'hxxxx;   // 193  -0.716  -0.698
    assign  wn_re[194] = 16'hA34C;   assign  wn_im[194] = 16'hA7BD;   // 194  -0.724  -0.690
    assign  wn_re[195] = 16'hA238;   assign  wn_im[195] = 16'hA8E2;   // 195  -0.733  -0.681
    assign  wn_re[196] = 16'hA129;   assign  wn_im[196] = 16'hAA0A;   // 196  -0.741  -0.672
    assign  wn_re[197] = 16'hxxxx;   assign  wn_im[197] = 16'hxxxx;   // 197  -0.749  -0.662
    assign  wn_re[198] = 16'h9F14;   assign  wn_im[198] = 16'hAC65;   // 198  -0.757  -0.653
    assign  wn_re[199] = 16'hxxxx;   assign  wn_im[199] = 16'hxxxx;   // 199  -0.765  -0.644
    assign  wn_re[200] = 16'h9D0E;   assign  wn_im[200] = 16'hAECC;   // 200  -0.773  -0.634
    assign  wn_re[201] = 16'h9C11;   assign  wn_im[201] = 16'hB005;   // 201  -0.781  -0.625
    assign  wn_re[202] = 16'h9B17;   assign  wn_im[202] = 16'hB140;   // 202  -0.788  -0.615
    assign  wn_re[203] = 16'hxxxx;   assign  wn_im[203] = 16'hxxxx;   // 203  -0.796  -0.606
    assign  wn_re[204] = 16'h9930;   assign  wn_im[204] = 16'hB3C0;   // 204  -0.803  -0.596
    assign  wn_re[205] = 16'hxxxx;   assign  wn_im[205] = 16'hxxxx;   // 205  -0.810  -0.586
    assign  wn_re[206] = 16'h9759;   assign  wn_im[206] = 16'hB64C;   // 206  -0.818  -0.576
    assign  wn_re[207] = 16'h9674;   assign  wn_im[207] = 16'hB796;   // 207  -0.825  -0.566
    assign  wn_re[208] = 16'h9592;   assign  wn_im[208] = 16'hB8E3;   // 208  -0.831  -0.556
    assign  wn_re[209] = 16'hxxxx;   assign  wn_im[209] = 16'hxxxx;   // 209  -0.838  -0.545
    assign  wn_re[210] = 16'h93DC;   assign  wn_im[210] = 16'hBB85;   // 210  -0.845  -0.535
    assign  wn_re[211] = 16'hxxxx;   assign  wn_im[211] = 16'hxxxx;   // 211  -0.851  -0.525
    assign  wn_re[212] = 16'h9236;   assign  wn_im[212] = 16'hBE32;   // 212  -0.858  -0.514
    assign  wn_re[213] = 16'h9169;   assign  wn_im[213] = 16'hBF8C;   // 213  -0.864  -0.504
    assign  wn_re[214] = 16'h90A1;   assign  wn_im[214] = 16'hC0E9;   // 214  -0.870  -0.493
    assign  wn_re[215] = 16'hxxxx;   assign  wn_im[215] = 16'hxxxx;   // 215  -0.876  -0.482
    assign  wn_re[216] = 16'h8F1D;   assign  wn_im[216] = 16'hC3A9;   // 216  -0.882  -0.471
    assign  wn_re[217] = 16'hxxxx;   assign  wn_im[217] = 16'hxxxx;   // 217  -0.888  -0.461
    assign  wn_re[218] = 16'h8DAB;   assign  wn_im[218] = 16'hC673;   // 218  -0.893  -0.450
    assign  wn_re[219] = 16'h8CF8;   assign  wn_im[219] = 16'hC7DB;   // 219  -0.899  -0.439
    assign  wn_re[220] = 16'h8C4A;   assign  wn_im[220] = 16'hC946;   // 220  -0.904  -0.428
    assign  wn_re[221] = 16'hxxxx;   assign  wn_im[221] = 16'hxxxx;   // 221  -0.909  -0.416
    assign  wn_re[222] = 16'h8AFB;   assign  wn_im[222] = 16'hCC21;   // 222  -0.914  -0.405
    assign  wn_re[223] = 16'hxxxx;   assign  wn_im[223] = 16'hxxxx;   // 223  -0.919  -0.394
    assign  wn_re[224] = 16'h89BE;   assign  wn_im[224] = 16'hCF04;   // 224  -0.924  -0.383
    assign  wn_re[225] = 16'h8927;   assign  wn_im[225] = 16'hD079;   // 225  -0.929  -0.371
    assign  wn_re[226] = 16'h8894;   assign  wn_im[226] = 16'hD1EF;   // 226  -0.933  -0.360
    assign  wn_re[227] = 16'hxxxx;   assign  wn_im[227] = 16'hxxxx;   // 227  -0.937  -0.348
    assign  wn_re[228] = 16'h877B;   assign  wn_im[228] = 16'hD4E1;   // 228  -0.942  -0.337
    assign  wn_re[229] = 16'hxxxx;   assign  wn_im[229] = 16'hxxxx;   // 229  -0.946  -0.325
    assign  wn_re[230] = 16'h8676;   assign  wn_im[230] = 16'hD7D9;   // 230  -0.950  -0.314
    assign  wn_re[231] = 16'h85FA;   assign  wn_im[231] = 16'hD958;   // 231  -0.953  -0.302
    assign  wn_re[232] = 16'h8583;   assign  wn_im[232] = 16'hDAD8;   // 232  -0.957  -0.290
    assign  wn_re[233] = 16'hxxxx;   assign  wn_im[233] = 16'hxxxx;   // 233  -0.960  -0.279
    assign  wn_re[234] = 16'h84A3;   assign  wn_im[234] = 16'hDDDC;   // 234  -0.964  -0.267
    assign  wn_re[235] = 16'hxxxx;   assign  wn_im[235] = 16'hxxxx;   // 235  -0.967  -0.255
    assign  wn_re[236] = 16'h83D6;   assign  wn_im[236] = 16'hE0E6;   // 236  -0.970  -0.243
    assign  wn_re[237] = 16'h8377;   assign  wn_im[237] = 16'hE26D;   // 237  -0.973  -0.231
    assign  wn_re[238] = 16'h831C;   assign  wn_im[238] = 16'hE3F4;   // 238  -0.976  -0.219
    assign  wn_re[239] = 16'hxxxx;   assign  wn_im[239] = 16'hxxxx;   // 239  -0.978  -0.207
    assign  wn_re[240] = 16'h8276;   assign  wn_im[240] = 16'hE707;   // 240  -0.981  -0.195
    assign  wn_re[241] = 16'hxxxx;   assign  wn_im[241] = 16'hxxxx;   // 241  -0.983  -0.183
    assign  wn_re[242] = 16'h81E2;   assign  wn_im[242] = 16'hEA1E;   // 242  -0.985  -0.171
    assign  wn_re[243] = 16'h81A0;   assign  wn_im[243] = 16'hEBAB;   // 243  -0.987  -0.159
    assign  wn_re[244] = 16'h8163;   assign  wn_im[244] = 16'hED38;   // 244  -0.989  -0.147
    assign  wn_re[245] = 16'hxxxx;   assign  wn_im[245] = 16'hxxxx;   // 245  -0.991  -0.135
    assign  wn_re[246] = 16'h80F6;   assign  wn_im[246] = 16'hF055;   // 246  -0.992  -0.122
    assign  wn_re[247] = 16'hxxxx;   assign  wn_im[247] = 16'hxxxx;   // 247  -0.994  -0.110
    assign  wn_re[248] = 16'h809E;   assign  wn_im[248] = 16'hF374;   // 248  -0.995  -0.098
    assign  wn_re[249] = 16'h8079;   assign  wn_im[249] = 16'hF505;   // 249  -0.996  -0.086
    assign  wn_re[250] = 16'h8059;   assign  wn_im[250] = 16'hF695;   // 250  -0.997  -0.074
    assign  wn_re[251] = 16'hxxxx;   assign  wn_im[251] = 16'hxxxx;   // 251  -0.998  -0.061
    assign  wn_re[252] = 16'h8027;   assign  wn_im[252] = 16'hF9B8;   // 252  -0.999  -0.049
    assign  wn_re[253] = 16'hxxxx;   assign  wn_im[253] = 16'hxxxx;   // 253  -0.999  -0.037
    assign  wn_re[254] = 16'h800A;   assign  wn_im[254] = 16'hFCDC;   // 254  -1.000  -0.025
    assign  wn_re[255] = 16'h8002;   assign  wn_im[255] = 16'hFE6E;   // 255  -1.000  -0.012
    assign  wn_re[256] = 16'hxxxx;   assign  wn_im[256] = 16'hxxxx;   // 256  -1.000  -0.000
    assign  wn_re[257] = 16'hxxxx;   assign  wn_im[257] = 16'hxxxx;   // 257  -1.000   0.012
    assign  wn_re[258] = 16'h800A;   assign  wn_im[258] = 16'h0324;   // 258  -1.000   0.025
    assign  wn_re[259] = 16'hxxxx;   assign  wn_im[259] = 16'hxxxx;   // 259  -0.999   0.037
    assign  wn_re[260] = 16'hxxxx;   assign  wn_im[260] = 16'hxxxx;   // 260  -0.999   0.049
    assign  wn_re[261] = 16'h803E;   assign  wn_im[261] = 16'h07D9;   // 261  -0.998   0.061
    assign  wn_re[262] = 16'hxxxx;   assign  wn_im[262] = 16'hxxxx;   // 262  -0.997   0.074
    assign  wn_re[263] = 16'hxxxx;   assign  wn_im[263] = 16'hxxxx;   // 263  -0.996   0.086
    assign  wn_re[264] = 16'h809E;   assign  wn_im[264] = 16'h0C8C;   // 264  -0.995   0.098
    assign  wn_re[265] = 16'hxxxx;   assign  wn_im[265] = 16'hxxxx;   // 265  -0.994   0.110
    assign  wn_re[266] = 16'hxxxx;   assign  wn_im[266] = 16'hxxxx;   // 266  -0.992   0.122
    assign  wn_re[267] = 16'h812A;   assign  wn_im[267] = 16'h113A;   // 267  -0.991   0.135
    assign  wn_re[268] = 16'hxxxx;   assign  wn_im[268] = 16'hxxxx;   // 268  -0.989   0.147
    assign  wn_re[269] = 16'hxxxx;   assign  wn_im[269] = 16'hxxxx;   // 269  -0.987   0.159
    assign  wn_re[270] = 16'h81E2;   assign  wn_im[270] = 16'h15E2;   // 270  -0.985   0.171
    assign  wn_re[271] = 16'hxxxx;   assign  wn_im[271] = 16'hxxxx;   // 271  -0.983   0.183
    assign  wn_re[272] = 16'hxxxx;   assign  wn_im[272] = 16'hxxxx;   // 272  -0.981   0.195
    assign  wn_re[273] = 16'h82C6;   assign  wn_im[273] = 16'h1A83;   // 273  -0.978   0.207
    assign  wn_re[274] = 16'hxxxx;   assign  wn_im[274] = 16'hxxxx;   // 274  -0.976   0.219
    assign  wn_re[275] = 16'hxxxx;   assign  wn_im[275] = 16'hxxxx;   // 275  -0.973   0.231
    assign  wn_re[276] = 16'h83D6;   assign  wn_im[276] = 16'h1F1A;   // 276  -0.970   0.243
    assign  wn_re[277] = 16'hxxxx;   assign  wn_im[277] = 16'hxxxx;   // 277  -0.967   0.255
    assign  wn_re[278] = 16'hxxxx;   assign  wn_im[278] = 16'hxxxx;   // 278  -0.964   0.267
    assign  wn_re[279] = 16'h8511;   assign  wn_im[279] = 16'h23A7;   // 279  -0.960   0.279
    assign  wn_re[280] = 16'hxxxx;   assign  wn_im[280] = 16'hxxxx;   // 280  -0.957   0.290
    assign  wn_re[281] = 16'hxxxx;   assign  wn_im[281] = 16'hxxxx;   // 281  -0.953   0.302
    assign  wn_re[282] = 16'h8676;   assign  wn_im[282] = 16'h2827;   // 282  -0.950   0.314
    assign  wn_re[283] = 16'hxxxx;   assign  wn_im[283] = 16'hxxxx;   // 283  -0.946   0.325
    assign  wn_re[284] = 16'hxxxx;   assign  wn_im[284] = 16'hxxxx;   // 284  -0.942   0.337
    assign  wn_re[285] = 16'h8805;   assign  wn_im[285] = 16'h2C99;   // 285  -0.937   0.348
    assign  wn_re[286] = 16'hxxxx;   assign  wn_im[286] = 16'hxxxx;   // 286  -0.933   0.360
    assign  wn_re[287] = 16'hxxxx;   assign  wn_im[287] = 16'hxxxx;   // 287  -0.929   0.371
    assign  wn_re[288] = 16'h89BE;   assign  wn_im[288] = 16'h30FC;   // 288  -0.924   0.383
    assign  wn_re[289] = 16'hxxxx;   assign  wn_im[289] = 16'hxxxx;   // 289  -0.919   0.394
    assign  wn_re[290] = 16'hxxxx;   assign  wn_im[290] = 16'hxxxx;   // 290  -0.914   0.405
    assign  wn_re[291] = 16'h8BA0;   assign  wn_im[291] = 16'h354E;   // 291  -0.909   0.416
    assign  wn_re[292] = 16'hxxxx;   assign  wn_im[292] = 16'hxxxx;   // 292  -0.904   0.428
    assign  wn_re[293] = 16'hxxxx;   assign  wn_im[293] = 16'hxxxx;   // 293  -0.899   0.439
    assign  wn_re[294] = 16'h8DAB;   assign  wn_im[294] = 16'h398D;   // 294  -0.893   0.450
    assign  wn_re[295] = 16'hxxxx;   assign  wn_im[295] = 16'hxxxx;   // 295  -0.888   0.461
    assign  wn_re[296] = 16'hxxxx;   assign  wn_im[296] = 16'hxxxx;   // 296  -0.882   0.471
    assign  wn_re[297] = 16'h8FDD;   assign  wn_im[297] = 16'h3DB8;   // 297  -0.876   0.482
    assign  wn_re[298] = 16'hxxxx;   assign  wn_im[298] = 16'hxxxx;   // 298  -0.870   0.493
    assign  wn_re[299] = 16'hxxxx;   assign  wn_im[299] = 16'hxxxx;   // 299  -0.864   0.504
    assign  wn_re[300] = 16'h9236;   assign  wn_im[300] = 16'h41CE;   // 300  -0.858   0.514
    assign  wn_re[301] = 16'hxxxx;   assign  wn_im[301] = 16'hxxxx;   // 301  -0.851   0.525
    assign  wn_re[302] = 16'hxxxx;   assign  wn_im[302] = 16'hxxxx;   // 302  -0.845   0.535
    assign  wn_re[303] = 16'h94B5;   assign  wn_im[303] = 16'h45CD;   // 303  -0.838   0.545
    assign  wn_re[304] = 16'hxxxx;   assign  wn_im[304] = 16'hxxxx;   // 304  -0.831   0.556
    assign  wn_re[305] = 16'hxxxx;   assign  wn_im[305] = 16'hxxxx;   // 305  -0.825   0.566
    assign  wn_re[306] = 16'h9759;   assign  wn_im[306] = 16'h49B4;   // 306  -0.818   0.576
    assign  wn_re[307] = 16'hxxxx;   assign  wn_im[307] = 16'hxxxx;   // 307  -0.810   0.586
    assign  wn_re[308] = 16'hxxxx;   assign  wn_im[308] = 16'hxxxx;   // 308  -0.803   0.596
    assign  wn_re[309] = 16'h9A22;   assign  wn_im[309] = 16'h4D81;   // 309  -0.796   0.606
    assign  wn_re[310] = 16'hxxxx;   assign  wn_im[310] = 16'hxxxx;   // 310  -0.788   0.615
    assign  wn_re[311] = 16'hxxxx;   assign  wn_im[311] = 16'hxxxx;   // 311  -0.781   0.625
    assign  wn_re[312] = 16'h9D0E;   assign  wn_im[312] = 16'h5134;   // 312  -0.773   0.634
    assign  wn_re[313] = 16'hxxxx;   assign  wn_im[313] = 16'hxxxx;   // 313  -0.765   0.644
    assign  wn_re[314] = 16'hxxxx;   assign  wn_im[314] = 16'hxxxx;   // 314  -0.757   0.653
    assign  wn_re[315] = 16'hA01C;   assign  wn_im[315] = 16'h54CA;   // 315  -0.749   0.662
    assign  wn_re[316] = 16'hxxxx;   assign  wn_im[316] = 16'hxxxx;   // 316  -0.741   0.672
    assign  wn_re[317] = 16'hxxxx;   assign  wn_im[317] = 16'hxxxx;   // 317  -0.733   0.681
    assign  wn_re[318] = 16'hA34C;   assign  wn_im[318] = 16'h5843;   // 318  -0.724   0.690
    assign  wn_re[319] = 16'hxxxx;   assign  wn_im[319] = 16'hxxxx;   // 319  -0.716   0.698
    assign  wn_re[320] = 16'hxxxx;   assign  wn_im[320] = 16'hxxxx;   // 320  -0.707   0.707
    assign  wn_re[321] = 16'hA69C;   assign  wn_im[321] = 16'h5B9D;   // 321  -0.698   0.716
    assign  wn_re[322] = 16'hxxxx;   assign  wn_im[322] = 16'hxxxx;   // 322  -0.690   0.724
    assign  wn_re[323] = 16'hxxxx;   assign  wn_im[323] = 16'hxxxx;   // 323  -0.681   0.733
    assign  wn_re[324] = 16'hAA0A;   assign  wn_im[324] = 16'h5ED7;   // 324  -0.672   0.741
    assign  wn_re[325] = 16'hxxxx;   assign  wn_im[325] = 16'hxxxx;   // 325  -0.662   0.749
    assign  wn_re[326] = 16'hxxxx;   assign  wn_im[326] = 16'hxxxx;   // 326  -0.653   0.757
    assign  wn_re[327] = 16'hAD97;   assign  wn_im[327] = 16'h61F1;   // 327  -0.644   0.765
    assign  wn_re[328] = 16'hxxxx;   assign  wn_im[328] = 16'hxxxx;   // 328  -0.634   0.773
    assign  wn_re[329] = 16'hxxxx;   assign  wn_im[329] = 16'hxxxx;   // 329  -0.625   0.781
    assign  wn_re[330] = 16'hB140;   assign  wn_im[330] = 16'h64E9;   // 330  -0.615   0.788
    assign  wn_re[331] = 16'hxxxx;   assign  wn_im[331] = 16'hxxxx;   // 331  -0.606   0.796
    assign  wn_re[332] = 16'hxxxx;   assign  wn_im[332] = 16'hxxxx;   // 332  -0.596   0.803
    assign  wn_re[333] = 16'hB505;   assign  wn_im[333] = 16'h67BD;   // 333  -0.586   0.810
    assign  wn_re[334] = 16'hxxxx;   assign  wn_im[334] = 16'hxxxx;   // 334  -0.576   0.818
    assign  wn_re[335] = 16'hxxxx;   assign  wn_im[335] = 16'hxxxx;   // 335  -0.566   0.825
    assign  wn_re[336] = 16'hB8E3;   assign  wn_im[336] = 16'h6A6E;   // 336  -0.556   0.831
    assign  wn_re[337] = 16'hxxxx;   assign  wn_im[337] = 16'hxxxx;   // 337  -0.545   0.838
    assign  wn_re[338] = 16'hxxxx;   assign  wn_im[338] = 16'hxxxx;   // 338  -0.535   0.845
    assign  wn_re[339] = 16'hBCDA;   assign  wn_im[339] = 16'h6CF9;   // 339  -0.525   0.851
    assign  wn_re[340] = 16'hxxxx;   assign  wn_im[340] = 16'hxxxx;   // 340  -0.514   0.858
    assign  wn_re[341] = 16'hxxxx;   assign  wn_im[341] = 16'hxxxx;   // 341  -0.504   0.864
    assign  wn_re[342] = 16'hC0E9;   assign  wn_im[342] = 16'h6F5F;   // 342  -0.493   0.870
    assign  wn_re[343] = 16'hxxxx;   assign  wn_im[343] = 16'hxxxx;   // 343  -0.482   0.876
    assign  wn_re[344] = 16'hxxxx;   assign  wn_im[344] = 16'hxxxx;   // 344  -0.471   0.882
    assign  wn_re[345] = 16'hC50D;   assign  wn_im[345] = 16'h719E;   // 345  -0.461   0.888
    assign  wn_re[346] = 16'hxxxx;   assign  wn_im[346] = 16'hxxxx;   // 346  -0.450   0.893
    assign  wn_re[347] = 16'hxxxx;   assign  wn_im[347] = 16'hxxxx;   // 347  -0.439   0.899
    assign  wn_re[348] = 16'hC946;   assign  wn_im[348] = 16'h73B6;   // 348  -0.428   0.904
    assign  wn_re[349] = 16'hxxxx;   assign  wn_im[349] = 16'hxxxx;   // 349  -0.416   0.909
    assign  wn_re[350] = 16'hxxxx;   assign  wn_im[350] = 16'hxxxx;   // 350  -0.405   0.914
    assign  wn_re[351] = 16'hCD92;   assign  wn_im[351] = 16'h75A6;   // 351  -0.394   0.919
    assign  wn_re[352] = 16'hxxxx;   assign  wn_im[352] = 16'hxxxx;   // 352  -0.383   0.924
    assign  wn_re[353] = 16'hxxxx;   assign  wn_im[353] = 16'hxxxx;   // 353  -0.371   0.929
    assign  wn_re[354] = 16'hD1EF;   assign  wn_im[354] = 16'h776C;   // 354  -0.360   0.933
    assign  wn_re[355] = 16'hxxxx;   assign  wn_im[355] = 16'hxxxx;   // 355  -0.348   0.937
    assign  wn_re[356] = 16'hxxxx;   assign  wn_im[356] = 16'hxxxx;   // 356  -0.337   0.942
    assign  wn_re[357] = 16'hD65C;   assign  wn_im[357] = 16'h790A;   // 357  -0.325   0.946
    assign  wn_re[358] = 16'hxxxx;   assign  wn_im[358] = 16'hxxxx;   // 358  -0.314   0.950
    assign  wn_re[359] = 16'hxxxx;   assign  wn_im[359] = 16'hxxxx;   // 359  -0.302   0.953
    assign  wn_re[360] = 16'hDAD8;   assign  wn_im[360] = 16'h7A7D;   // 360  -0.290   0.957
    assign  wn_re[361] = 16'hxxxx;   assign  wn_im[361] = 16'hxxxx;   // 361  -0.279   0.960
    assign  wn_re[362] = 16'hxxxx;   assign  wn_im[362] = 16'hxxxx;   // 362  -0.267   0.964
    assign  wn_re[363] = 16'hDF61;   assign  wn_im[363] = 16'h7BC6;   // 363  -0.255   0.967
    assign  wn_re[364] = 16'hxxxx;   assign  wn_im[364] = 16'hxxxx;   // 364  -0.243   0.970
    assign  wn_re[365] = 16'hxxxx;   assign  wn_im[365] = 16'hxxxx;   // 365  -0.231   0.973
    assign  wn_re[366] = 16'hE3F4;   assign  wn_im[366] = 16'h7CE4;   // 366  -0.219   0.976
    assign  wn_re[367] = 16'hxxxx;   assign  wn_im[367] = 16'hxxxx;   // 367  -0.207   0.978
    assign  wn_re[368] = 16'hxxxx;   assign  wn_im[368] = 16'hxxxx;   // 368  -0.195   0.981
    assign  wn_re[369] = 16'hE892;   assign  wn_im[369] = 16'h7DD6;   // 369  -0.183   0.983
    assign  wn_re[370] = 16'hxxxx;   assign  wn_im[370] = 16'hxxxx;   // 370  -0.171   0.985
    assign  wn_re[371] = 16'hxxxx;   assign  wn_im[371] = 16'hxxxx;   // 371  -0.159   0.987
    assign  wn_re[372] = 16'hED38;   assign  wn_im[372] = 16'h7E9D;   // 372  -0.147   0.989
    assign  wn_re[373] = 16'hxxxx;   assign  wn_im[373] = 16'hxxxx;   // 373  -0.135   0.991
    assign  wn_re[374] = 16'hxxxx;   assign  wn_im[374] = 16'hxxxx;   // 374  -0.122   0.992
    assign  wn_re[375] = 16'hF1E4;   assign  wn_im[375] = 16'h7F38;   // 375  -0.110   0.994
    assign  wn_re[376] = 16'hxxxx;   assign  wn_im[376] = 16'hxxxx;   // 376  -0.098   0.995
    assign  wn_re[377] = 16'hxxxx;   assign  wn_im[377] = 16'hxxxx;   // 377  -0.086   0.996
    assign  wn_re[378] = 16'hF695;   assign  wn_im[378] = 16'h7FA7;   // 378  -0.074   0.997
    assign  wn_re[379] = 16'hxxxx;   assign  wn_im[379] = 16'hxxxx;   // 379  -0.061   0.998
    assign  wn_re[380] = 16'hxxxx;   assign  wn_im[380] = 16'hxxxx;   // 380  -0.049   0.999
    assign  wn_re[381] = 16'hFB4A;   assign  wn_im[381] = 16'h7FEA;   // 381  -0.037   0.999
    assign  wn_re[382] = 16'hxxxx;   assign  wn_im[382] = 16'hxxxx;   // 382  -0.025   1.000
    assign  wn_re[383] = 16'hxxxx;   assign  wn_im[383] = 16'hxxxx;   // 383  -0.012   1.000
    assign  wn_re[384] = 16'hxxxx;   assign  wn_im[384] = 16'hxxxx;   // 384  -0.000   1.000
    assign  wn_re[385] = 16'hxxxx;   assign  wn_im[385] = 16'hxxxx;   // 385   0.012   1.000
    assign  wn_re[386] = 16'hxxxx;   assign  wn_im[386] = 16'hxxxx;   // 386   0.025   1.000
    assign  wn_re[387] = 16'hxxxx;   assign  wn_im[387] = 16'hxxxx;   // 387   0.037   0.999
    assign  wn_re[388] = 16'hxxxx;   assign  wn_im[388] = 16'hxxxx;   // 388   0.049   0.999
    assign  wn_re[389] = 16'hxxxx;   assign  wn_im[389] = 16'hxxxx;   // 389   0.061   0.998
    assign  wn_re[390] = 16'hxxxx;   assign  wn_im[390] = 16'hxxxx;   // 390   0.074   0.997
    assign  wn_re[391] = 16'hxxxx;   assign  wn_im[391] = 16'hxxxx;   // 391   0.086   0.996
    assign  wn_re[392] = 16'hxxxx;   assign  wn_im[392] = 16'hxxxx;   // 392   0.098   0.995
    assign  wn_re[393] = 16'hxxxx;   assign  wn_im[393] = 16'hxxxx;   // 393   0.110   0.994
    assign  wn_re[394] = 16'hxxxx;   assign  wn_im[394] = 16'hxxxx;   // 394   0.122   0.992
    assign  wn_re[395] = 16'hxxxx;   assign  wn_im[395] = 16'hxxxx;   // 395   0.135   0.991
    assign  wn_re[396] = 16'hxxxx;   assign  wn_im[396] = 16'hxxxx;   // 396   0.147   0.989
    assign  wn_re[397] = 16'hxxxx;   assign  wn_im[397] = 16'hxxxx;   // 397   0.159   0.987
    assign  wn_re[398] = 16'hxxxx;   assign  wn_im[398] = 16'hxxxx;   // 398   0.171   0.985
    assign  wn_re[399] = 16'hxxxx;   assign  wn_im[399] = 16'hxxxx;   // 399   0.183   0.983
    assign  wn_re[400] = 16'hxxxx;   assign  wn_im[400] = 16'hxxxx;   // 400   0.195   0.981
    assign  wn_re[401] = 16'hxxxx;   assign  wn_im[401] = 16'hxxxx;   // 401   0.207   0.978
    assign  wn_re[402] = 16'hxxxx;   assign  wn_im[402] = 16'hxxxx;   // 402   0.219   0.976
    assign  wn_re[403] = 16'hxxxx;   assign  wn_im[403] = 16'hxxxx;   // 403   0.231   0.973
    assign  wn_re[404] = 16'hxxxx;   assign  wn_im[404] = 16'hxxxx;   // 404   0.243   0.970
    assign  wn_re[405] = 16'hxxxx;   assign  wn_im[405] = 16'hxxxx;   // 405   0.255   0.967
    assign  wn_re[406] = 16'hxxxx;   assign  wn_im[406] = 16'hxxxx;   // 406   0.267   0.964
    assign  wn_re[407] = 16'hxxxx;   assign  wn_im[407] = 16'hxxxx;   // 407   0.279   0.960
    assign  wn_re[408] = 16'hxxxx;   assign  wn_im[408] = 16'hxxxx;   // 408   0.290   0.957
    assign  wn_re[409] = 16'hxxxx;   assign  wn_im[409] = 16'hxxxx;   // 409   0.302   0.953
    assign  wn_re[410] = 16'hxxxx;   assign  wn_im[410] = 16'hxxxx;   // 410   0.314   0.950
    assign  wn_re[411] = 16'hxxxx;   assign  wn_im[411] = 16'hxxxx;   // 411   0.325   0.946
    assign  wn_re[412] = 16'hxxxx;   assign  wn_im[412] = 16'hxxxx;   // 412   0.337   0.942
    assign  wn_re[413] = 16'hxxxx;   assign  wn_im[413] = 16'hxxxx;   // 413   0.348   0.937
    assign  wn_re[414] = 16'hxxxx;   assign  wn_im[414] = 16'hxxxx;   // 414   0.360   0.933
    assign  wn_re[415] = 16'hxxxx;   assign  wn_im[415] = 16'hxxxx;   // 415   0.371   0.929
    assign  wn_re[416] = 16'hxxxx;   assign  wn_im[416] = 16'hxxxx;   // 416   0.383   0.924
    assign  wn_re[417] = 16'hxxxx;   assign  wn_im[417] = 16'hxxxx;   // 417   0.394   0.919
    assign  wn_re[418] = 16'hxxxx;   assign  wn_im[418] = 16'hxxxx;   // 418   0.405   0.914
    assign  wn_re[419] = 16'hxxxx;   assign  wn_im[419] = 16'hxxxx;   // 419   0.416   0.909
    assign  wn_re[420] = 16'hxxxx;   assign  wn_im[420] = 16'hxxxx;   // 420   0.428   0.904
    assign  wn_re[421] = 16'hxxxx;   assign  wn_im[421] = 16'hxxxx;   // 421   0.439   0.899
    assign  wn_re[422] = 16'hxxxx;   assign  wn_im[422] = 16'hxxxx;   // 422   0.450   0.893
    assign  wn_re[423] = 16'hxxxx;   assign  wn_im[423] = 16'hxxxx;   // 423   0.461   0.888
    assign  wn_re[424] = 16'hxxxx;   assign  wn_im[424] = 16'hxxxx;   // 424   0.471   0.882
    assign  wn_re[425] = 16'hxxxx;   assign  wn_im[425] = 16'hxxxx;   // 425   0.482   0.876
    assign  wn_re[426] = 16'hxxxx;   assign  wn_im[426] = 16'hxxxx;   // 426   0.493   0.870
    assign  wn_re[427] = 16'hxxxx;   assign  wn_im[427] = 16'hxxxx;   // 427   0.504   0.864
    assign  wn_re[428] = 16'hxxxx;   assign  wn_im[428] = 16'hxxxx;   // 428   0.514   0.858
    assign  wn_re[429] = 16'hxxxx;   assign  wn_im[429] = 16'hxxxx;   // 429   0.525   0.851
    assign  wn_re[430] = 16'hxxxx;   assign  wn_im[430] = 16'hxxxx;   // 430   0.535   0.845
    assign  wn_re[431] = 16'hxxxx;   assign  wn_im[431] = 16'hxxxx;   // 431   0.545   0.838
    assign  wn_re[432] = 16'hxxxx;   assign  wn_im[432] = 16'hxxxx;   // 432   0.556   0.831
    assign  wn_re[433] = 16'hxxxx;   assign  wn_im[433] = 16'hxxxx;   // 433   0.566   0.825
    assign  wn_re[434] = 16'hxxxx;   assign  wn_im[434] = 16'hxxxx;   // 434   0.576   0.818
    assign  wn_re[435] = 16'hxxxx;   assign  wn_im[435] = 16'hxxxx;   // 435   0.586   0.810
    assign  wn_re[436] = 16'hxxxx;   assign  wn_im[436] = 16'hxxxx;   // 436   0.596   0.803
    assign  wn_re[437] = 16'hxxxx;   assign  wn_im[437] = 16'hxxxx;   // 437   0.606   0.796
    assign  wn_re[438] = 16'hxxxx;   assign  wn_im[438] = 16'hxxxx;   // 438   0.615   0.788
    assign  wn_re[439] = 16'hxxxx;   assign  wn_im[439] = 16'hxxxx;   // 439   0.625   0.781
    assign  wn_re[440] = 16'hxxxx;   assign  wn_im[440] = 16'hxxxx;   // 440   0.634   0.773
    assign  wn_re[441] = 16'hxxxx;   assign  wn_im[441] = 16'hxxxx;   // 441   0.644   0.765
    assign  wn_re[442] = 16'hxxxx;   assign  wn_im[442] = 16'hxxxx;   // 442   0.653   0.757
    assign  wn_re[443] = 16'hxxxx;   assign  wn_im[443] = 16'hxxxx;   // 443   0.662   0.749
    assign  wn_re[444] = 16'hxxxx;   assign  wn_im[444] = 16'hxxxx;   // 444   0.672   0.741
    assign  wn_re[445] = 16'hxxxx;   assign  wn_im[445] = 16'hxxxx;   // 445   0.681   0.733
    assign  wn_re[446] = 16'hxxxx;   assign  wn_im[446] = 16'hxxxx;   // 446   0.690   0.724
    assign  wn_re[447] = 16'hxxxx;   assign  wn_im[447] = 16'hxxxx;   // 447   0.698   0.716
    assign  wn_re[448] = 16'hxxxx;   assign  wn_im[448] = 16'hxxxx;   // 448   0.707   0.707
    assign  wn_re[449] = 16'hxxxx;   assign  wn_im[449] = 16'hxxxx;   // 449   0.716   0.698
    assign  wn_re[450] = 16'hxxxx;   assign  wn_im[450] = 16'hxxxx;   // 450   0.724   0.690
    assign  wn_re[451] = 16'hxxxx;   assign  wn_im[451] = 16'hxxxx;   // 451   0.733   0.681
    assign  wn_re[452] = 16'hxxxx;   assign  wn_im[452] = 16'hxxxx;   // 452   0.741   0.672
    assign  wn_re[453] = 16'hxxxx;   assign  wn_im[453] = 16'hxxxx;   // 453   0.749   0.662
    assign  wn_re[454] = 16'hxxxx;   assign  wn_im[454] = 16'hxxxx;   // 454   0.757   0.653
    assign  wn_re[455] = 16'hxxxx;   assign  wn_im[455] = 16'hxxxx;   // 455   0.765   0.644
    assign  wn_re[456] = 16'hxxxx;   assign  wn_im[456] = 16'hxxxx;   // 456   0.773   0.634
    assign  wn_re[457] = 16'hxxxx;   assign  wn_im[457] = 16'hxxxx;   // 457   0.781   0.625
    assign  wn_re[458] = 16'hxxxx;   assign  wn_im[458] = 16'hxxxx;   // 458   0.788   0.615
    assign  wn_re[459] = 16'hxxxx;   assign  wn_im[459] = 16'hxxxx;   // 459   0.796   0.606
    assign  wn_re[460] = 16'hxxxx;   assign  wn_im[460] = 16'hxxxx;   // 460   0.803   0.596
    assign  wn_re[461] = 16'hxxxx;   assign  wn_im[461] = 16'hxxxx;   // 461   0.810   0.586
    assign  wn_re[462] = 16'hxxxx;   assign  wn_im[462] = 16'hxxxx;   // 462   0.818   0.576
    assign  wn_re[463] = 16'hxxxx;   assign  wn_im[463] = 16'hxxxx;   // 463   0.825   0.566
    assign  wn_re[464] = 16'hxxxx;   assign  wn_im[464] = 16'hxxxx;   // 464   0.831   0.556
    assign  wn_re[465] = 16'hxxxx;   assign  wn_im[465] = 16'hxxxx;   // 465   0.838   0.545
    assign  wn_re[466] = 16'hxxxx;   assign  wn_im[466] = 16'hxxxx;   // 466   0.845   0.535
    assign  wn_re[467] = 16'hxxxx;   assign  wn_im[467] = 16'hxxxx;   // 467   0.851   0.525
    assign  wn_re[468] = 16'hxxxx;   assign  wn_im[468] = 16'hxxxx;   // 468   0.858   0.514
    assign  wn_re[469] = 16'hxxxx;   assign  wn_im[469] = 16'hxxxx;   // 469   0.864   0.504
    assign  wn_re[470] = 16'hxxxx;   assign  wn_im[470] = 16'hxxxx;   // 470   0.870   0.493
    assign  wn_re[471] = 16'hxxxx;   assign  wn_im[471] = 16'hxxxx;   // 471   0.876   0.482
    assign  wn_re[472] = 16'hxxxx;   assign  wn_im[472] = 16'hxxxx;   // 472   0.882   0.471
    assign  wn_re[473] = 16'hxxxx;   assign  wn_im[473] = 16'hxxxx;   // 473   0.888   0.461
    assign  wn_re[474] = 16'hxxxx;   assign  wn_im[474] = 16'hxxxx;   // 474   0.893   0.450
    assign  wn_re[475] = 16'hxxxx;   assign  wn_im[475] = 16'hxxxx;   // 475   0.899   0.439
    assign  wn_re[476] = 16'hxxxx;   assign  wn_im[476] = 16'hxxxx;   // 476   0.904   0.428
    assign  wn_re[477] = 16'hxxxx;   assign  wn_im[477] = 16'hxxxx;   // 477   0.909   0.416
    assign  wn_re[478] = 16'hxxxx;   assign  wn_im[478] = 16'hxxxx;   // 478   0.914   0.405
    assign  wn_re[479] = 16'hxxxx;   assign  wn_im[479] = 16'hxxxx;   // 479   0.919   0.394
    assign  wn_re[480] = 16'hxxxx;   assign  wn_im[480] = 16'hxxxx;   // 480   0.924   0.383
    assign  wn_re[481] = 16'hxxxx;   assign  wn_im[481] = 16'hxxxx;   // 481   0.929   0.371
    assign  wn_re[482] = 16'hxxxx;   assign  wn_im[482] = 16'hxxxx;   // 482   0.933   0.360
    assign  wn_re[483] = 16'hxxxx;   assign  wn_im[483] = 16'hxxxx;   // 483   0.937   0.348
    assign  wn_re[484] = 16'hxxxx;   assign  wn_im[484] = 16'hxxxx;   // 484   0.942   0.337
    assign  wn_re[485] = 16'hxxxx;   assign  wn_im[485] = 16'hxxxx;   // 485   0.946   0.325
    assign  wn_re[486] = 16'hxxxx;   assign  wn_im[486] = 16'hxxxx;   // 486   0.950   0.314
    assign  wn_re[487] = 16'hxxxx;   assign  wn_im[487] = 16'hxxxx;   // 487   0.953   0.302
    assign  wn_re[488] = 16'hxxxx;   assign  wn_im[488] = 16'hxxxx;   // 488   0.957   0.290
    assign  wn_re[489] = 16'hxxxx;   assign  wn_im[489] = 16'hxxxx;   // 489   0.960   0.279
    assign  wn_re[490] = 16'hxxxx;   assign  wn_im[490] = 16'hxxxx;   // 490   0.964   0.267
    assign  wn_re[491] = 16'hxxxx;   assign  wn_im[491] = 16'hxxxx;   // 491   0.967   0.255
    assign  wn_re[492] = 16'hxxxx;   assign  wn_im[492] = 16'hxxxx;   // 492   0.970   0.243
    assign  wn_re[493] = 16'hxxxx;   assign  wn_im[493] = 16'hxxxx;   // 493   0.973   0.231
    assign  wn_re[494] = 16'hxxxx;   assign  wn_im[494] = 16'hxxxx;   // 494   0.976   0.219
    assign  wn_re[495] = 16'hxxxx;   assign  wn_im[495] = 16'hxxxx;   // 495   0.978   0.207
    assign  wn_re[496] = 16'hxxxx;   assign  wn_im[496] = 16'hxxxx;   // 496   0.981   0.195
    assign  wn_re[497] = 16'hxxxx;   assign  wn_im[497] = 16'hxxxx;   // 497   0.983   0.183
    assign  wn_re[498] = 16'hxxxx;   assign  wn_im[498] = 16'hxxxx;   // 498   0.985   0.171
    assign  wn_re[499] = 16'hxxxx;   assign  wn_im[499] = 16'hxxxx;   // 499   0.987   0.159
    assign  wn_re[500] = 16'hxxxx;   assign  wn_im[500] = 16'hxxxx;   // 500   0.989   0.147
    assign  wn_re[501] = 16'hxxxx;   assign  wn_im[501] = 16'hxxxx;   // 501   0.991   0.135
    assign  wn_re[502] = 16'hxxxx;   assign  wn_im[502] = 16'hxxxx;   // 502   0.992   0.122
    assign  wn_re[503] = 16'hxxxx;   assign  wn_im[503] = 16'hxxxx;   // 503   0.994   0.110
    assign  wn_re[504] = 16'hxxxx;   assign  wn_im[504] = 16'hxxxx;   // 504   0.995   0.098
    assign  wn_re[505] = 16'hxxxx;   assign  wn_im[505] = 16'hxxxx;   // 505   0.996   0.086
    assign  wn_re[506] = 16'hxxxx;   assign  wn_im[506] = 16'hxxxx;   // 506   0.997   0.074
    assign  wn_re[507] = 16'hxxxx;   assign  wn_im[507] = 16'hxxxx;   // 507   0.998   0.061
    assign  wn_re[508] = 16'hxxxx;   assign  wn_im[508] = 16'hxxxx;   // 508   0.999   0.049
    assign  wn_re[509] = 16'hxxxx;   assign  wn_im[509] = 16'hxxxx;   // 509   0.999   0.037
    assign  wn_re[510] = 16'hxxxx;   assign  wn_im[510] = 16'hxxxx;   // 510   1.000   0.025
    assign  wn_re[511] = 16'hxxxx;   assign  wn_im[511] = 16'hxxxx;   // 511   1.000   0.012

endmodule