// Hann Window Coefficients
// Length: 512
// Bit Width: 16
// Max Value: 32767
module HANN_WIN_480#(
    parameter N_FFT        = 512,
    parameter WIN_LEN      = 480,
    parameter ADDR_WIDTH = $clog2(N_FFT)
)( 
    input                   clk,
    input                   rst_n,
    input [ADDR_WIDTH-1:0]  addr,
    output reg [15:0]       win_coe_out
);

    

    
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            win_coe_out <= 16'h0000;
        end else begin
            win_coe_out <= addr < WIN_LEN ? win_coe[addr] : 16'h0000;
        end 
    end 
    
    wire [15:0] win_coe [0:N_FFT-1];

    assign win_coe [  0] = 16'h0000;
    assign win_coe [  1] = 16'h0001;
    assign win_coe [  2] = 16'h0006;
    assign win_coe [  3] = 16'h000d;
    assign win_coe [  4] = 16'h0017;
    assign win_coe [  5] = 16'h0023;
    assign win_coe [  6] = 16'h0033;
    assign win_coe [  7] = 16'h0045;
    assign win_coe [  8] = 16'h005a;
    assign win_coe [  9] = 16'h0072;
    assign win_coe [ 10] = 16'h008d;
    assign win_coe [ 11] = 16'h00aa;
    assign win_coe [ 12] = 16'h00cb;
    assign win_coe [ 13] = 16'h00ee;
    assign win_coe [ 14] = 16'h0113;
    assign win_coe [ 15] = 16'h013c;
    assign win_coe [ 16] = 16'h0168;
    assign win_coe [ 17] = 16'h0196;
    assign win_coe [ 18] = 16'h01c7;
    assign win_coe [ 19] = 16'h01fa;
    assign win_coe [ 20] = 16'h0231;
    assign win_coe [ 21] = 16'h026a;
    assign win_coe [ 22] = 16'h02a5;
    assign win_coe [ 23] = 16'h02e4;
    assign win_coe [ 24] = 16'h0325;
    assign win_coe [ 25] = 16'h0369;
    assign win_coe [ 26] = 16'h03b0;
    assign win_coe [ 27] = 16'h03f9;
    assign win_coe [ 28] = 16'h0445;
    assign win_coe [ 29] = 16'h0493;
    assign win_coe [ 30] = 16'h04e4;
    assign win_coe [ 31] = 16'h0538;
    assign win_coe [ 32] = 16'h058e;
    assign win_coe [ 33] = 16'h05e7;
    assign win_coe [ 34] = 16'h0643;
    assign win_coe [ 35] = 16'h06a1;
    assign win_coe [ 36] = 16'h0701;
    assign win_coe [ 37] = 16'h0764;
    assign win_coe [ 38] = 16'h07ca;
    assign win_coe [ 39] = 16'h0832;
    assign win_coe [ 40] = 16'h089c;
    assign win_coe [ 41] = 16'h0909;
    assign win_coe [ 42] = 16'h0978;
    assign win_coe [ 43] = 16'h09ea;
    assign win_coe [ 44] = 16'h0a5e;
    assign win_coe [ 45] = 16'h0ad4;
    assign win_coe [ 46] = 16'h0b4d;
    assign win_coe [ 47] = 16'h0bc8;
    assign win_coe [ 48] = 16'h0c46;
    assign win_coe [ 49] = 16'h0cc5;
    assign win_coe [ 50] = 16'h0d47;
    assign win_coe [ 51] = 16'h0dcb;
    assign win_coe [ 52] = 16'h0e52;
    assign win_coe [ 53] = 16'h0eda;
    assign win_coe [ 54] = 16'h0f65;
    assign win_coe [ 55] = 16'h0ff2;
    assign win_coe [ 56] = 16'h1081;
    assign win_coe [ 57] = 16'h1112;
    assign win_coe [ 58] = 16'h11a5;
    assign win_coe [ 59] = 16'h123a;
    assign win_coe [ 60] = 16'h12d2;
    assign win_coe [ 61] = 16'h136b;
    assign win_coe [ 62] = 16'h1406;
    assign win_coe [ 63] = 16'h14a3;
    assign win_coe [ 64] = 16'h1542;
    assign win_coe [ 65] = 16'h15e3;
    assign win_coe [ 66] = 16'h1686;
    assign win_coe [ 67] = 16'h172a;
    assign win_coe [ 68] = 16'h17d1;
    assign win_coe [ 69] = 16'h1879;
    assign win_coe [ 70] = 16'h1923;
    assign win_coe [ 71] = 16'h19ce;
    assign win_coe [ 72] = 16'h1a7c;
    assign win_coe [ 73] = 16'h1b2b;
    assign win_coe [ 74] = 16'h1bdb;
    assign win_coe [ 75] = 16'h1c8d;
    assign win_coe [ 76] = 16'h1d41;
    assign win_coe [ 77] = 16'h1df6;
    assign win_coe [ 78] = 16'h1ead;
    assign win_coe [ 79] = 16'h1f65;
    assign win_coe [ 80] = 16'h201f;
    assign win_coe [ 81] = 16'h20da;
    assign win_coe [ 82] = 16'h2196;
    assign win_coe [ 83] = 16'h2254;
    assign win_coe [ 84] = 16'h2313;
    assign win_coe [ 85] = 16'h23d3;
    assign win_coe [ 86] = 16'h2495;
    assign win_coe [ 87] = 16'h2558;
    assign win_coe [ 88] = 16'h261c;
    assign win_coe [ 89] = 16'h26e1;
    assign win_coe [ 90] = 16'h27a7;
    assign win_coe [ 91] = 16'h286e;
    assign win_coe [ 92] = 16'h2937;
    assign win_coe [ 93] = 16'h2a00;
    assign win_coe [ 94] = 16'h2aca;
    assign win_coe [ 95] = 16'h2b95;
    assign win_coe [ 96] = 16'h2c62;
    assign win_coe [ 97] = 16'h2d2f;
    assign win_coe [ 98] = 16'h2dfc;
    assign win_coe [ 99] = 16'h2ecb;
    assign win_coe [100] = 16'h2f9a;
    assign win_coe [101] = 16'h306a;
    assign win_coe [102] = 16'h313b;
    assign win_coe [103] = 16'h320d;
    assign win_coe [104] = 16'h32df;
    assign win_coe [105] = 16'h33b1;
    assign win_coe [106] = 16'h3485;
    assign win_coe [107] = 16'h3558;
    assign win_coe [108] = 16'h362c;
    assign win_coe [109] = 16'h3701;
    assign win_coe [110] = 16'h37d6;
    assign win_coe [111] = 16'h38ab;
    assign win_coe [112] = 16'h3981;
    assign win_coe [113] = 16'h3a57;
    assign win_coe [114] = 16'h3b2d;
    assign win_coe [115] = 16'h3c03;
    assign win_coe [116] = 16'h3cda;
    assign win_coe [117] = 16'h3db1;
    assign win_coe [118] = 16'h3e87;
    assign win_coe [119] = 16'h3f5e;
    assign win_coe [120] = 16'h4035;
    assign win_coe [121] = 16'h410c;
    assign win_coe [122] = 16'h41e3;
    assign win_coe [123] = 16'h42ba;
    assign win_coe [124] = 16'h4390;
    assign win_coe [125] = 16'h4467;
    assign win_coe [126] = 16'h453d;
    assign win_coe [127] = 16'h4613;
    assign win_coe [128] = 16'h46e9;
    assign win_coe [129] = 16'h47bf;
    assign win_coe [130] = 16'h4894;
    assign win_coe [131] = 16'h4968;
    assign win_coe [132] = 16'h4a3d;
    assign win_coe [133] = 16'h4b11;
    assign win_coe [134] = 16'h4be4;
    assign win_coe [135] = 16'h4cb7;
    assign win_coe [136] = 16'h4d89;
    assign win_coe [137] = 16'h4e5b;
    assign win_coe [138] = 16'h4f2c;
    assign win_coe [139] = 16'h4ffd;
    assign win_coe [140] = 16'h50cc;
    assign win_coe [141] = 16'h519b;
    assign win_coe [142] = 16'h526a;
    assign win_coe [143] = 16'h5337;
    assign win_coe [144] = 16'h5404;
    assign win_coe [145] = 16'h54cf;
    assign win_coe [146] = 16'h559a;
    assign win_coe [147] = 16'h5664;
    assign win_coe [148] = 16'h572d;
    assign win_coe [149] = 16'h57f4;
    assign win_coe [150] = 16'h58bb;
    assign win_coe [151] = 16'h5981;
    assign win_coe [152] = 16'h5a45;
    assign win_coe [153] = 16'h5b09;
    assign win_coe [154] = 16'h5bcb;
    assign win_coe [155] = 16'h5c8c;
    assign win_coe [156] = 16'h5d4c;
    assign win_coe [157] = 16'h5e0a;
    assign win_coe [158] = 16'h5ec7;
    assign win_coe [159] = 16'h5f83;
    assign win_coe [160] = 16'h603d;
    assign win_coe [161] = 16'h60f6;
    assign win_coe [162] = 16'h61ae;
    assign win_coe [163] = 16'h6264;
    assign win_coe [164] = 16'h6318;
    assign win_coe [165] = 16'h63cb;
    assign win_coe [166] = 16'h647c;
    assign win_coe [167] = 16'h652c;
    assign win_coe [168] = 16'h65da;
    assign win_coe [169] = 16'h6687;
    assign win_coe [170] = 16'h6731;
    assign win_coe [171] = 16'h67da;
    assign win_coe [172] = 16'h6882;
    assign win_coe [173] = 16'h6927;
    assign win_coe [174] = 16'h69cb;
    assign win_coe [175] = 16'h6a6d;
    assign win_coe [176] = 16'h6b0d;
    assign win_coe [177] = 16'h6bab;
    assign win_coe [178] = 16'h6c47;
    assign win_coe [179] = 16'h6ce1;
    assign win_coe [180] = 16'h6d79;
    assign win_coe [181] = 16'h6e0f;
    assign win_coe [182] = 16'h6ea4;
    assign win_coe [183] = 16'h6f36;
    assign win_coe [184] = 16'h6fc6;
    assign win_coe [185] = 16'h7054;
    assign win_coe [186] = 16'h70e0;
    assign win_coe [187] = 16'h7169;
    assign win_coe [188] = 16'h71f1;
    assign win_coe [189] = 16'h7276;
    assign win_coe [190] = 16'h72f9;
    assign win_coe [191] = 16'h737a;
    assign win_coe [192] = 16'h73f8;
    assign win_coe [193] = 16'h7475;
    assign win_coe [194] = 16'h74ef;
    assign win_coe [195] = 16'h7566;
    assign win_coe [196] = 16'h75db;
    assign win_coe [197] = 16'h764e;
    assign win_coe [198] = 16'h76bf;
    assign win_coe [199] = 16'h772d;
    assign win_coe [200] = 16'h7799;
    assign win_coe [201] = 16'h7802;
    assign win_coe [202] = 16'h7869;
    assign win_coe [203] = 16'h78cd;
    assign win_coe [204] = 16'h792f;
    assign win_coe [205] = 16'h798e;
    assign win_coe [206] = 16'h79ea;
    assign win_coe [207] = 16'h7a45;
    assign win_coe [208] = 16'h7a9c;
    assign win_coe [209] = 16'h7af1;
    assign win_coe [210] = 16'h7b44;
    assign win_coe [211] = 16'h7b93;
    assign win_coe [212] = 16'h7be1;
    assign win_coe [213] = 16'h7c2b;
    assign win_coe [214] = 16'h7c73;
    assign win_coe [215] = 16'h7cb8;
    assign win_coe [216] = 16'h7cfb;
    assign win_coe [217] = 16'h7d3b;
    assign win_coe [218] = 16'h7d78;
    assign win_coe [219] = 16'h7db2;
    assign win_coe [220] = 16'h7dea;
    assign win_coe [221] = 16'h7e1f;
    assign win_coe [222] = 16'h7e51;
    assign win_coe [223] = 16'h7e81;
    assign win_coe [224] = 16'h7eae;
    assign win_coe [225] = 16'h7ed8;
    assign win_coe [226] = 16'h7eff;
    assign win_coe [227] = 16'h7f23;
    assign win_coe [228] = 16'h7f45;
    assign win_coe [229] = 16'h7f64;
    assign win_coe [230] = 16'h7f80;
    assign win_coe [231] = 16'h7f99;
    assign win_coe [232] = 16'h7fb0;
    assign win_coe [233] = 16'h7fc3;
    assign win_coe [234] = 16'h7fd4;
    assign win_coe [235] = 16'h7fe2;
    assign win_coe [236] = 16'h7fee;
    assign win_coe [237] = 16'h7ff6;
    assign win_coe [238] = 16'h7ffc;
    assign win_coe [239] = 16'h7fff;
    assign win_coe [240] = 16'h7fff;
    assign win_coe [241] = 16'h7ffc;
    assign win_coe [242] = 16'h7ff6;
    assign win_coe [243] = 16'h7fee;
    assign win_coe [244] = 16'h7fe2;
    assign win_coe [245] = 16'h7fd4;
    assign win_coe [246] = 16'h7fc3;
    assign win_coe [247] = 16'h7fb0;
    assign win_coe [248] = 16'h7f99;
    assign win_coe [249] = 16'h7f80;
    assign win_coe [250] = 16'h7f64;
    assign win_coe [251] = 16'h7f45;
    assign win_coe [252] = 16'h7f23;
    assign win_coe [253] = 16'h7eff;
    assign win_coe [254] = 16'h7ed8;
    assign win_coe [255] = 16'h7eae;
    assign win_coe [256] = 16'h7e81;
    assign win_coe [257] = 16'h7e51;
    assign win_coe [258] = 16'h7e1f;
    assign win_coe [259] = 16'h7dea;
    assign win_coe [260] = 16'h7db2;
    assign win_coe [261] = 16'h7d78;
    assign win_coe [262] = 16'h7d3b;
    assign win_coe [263] = 16'h7cfb;
    assign win_coe [264] = 16'h7cb8;
    assign win_coe [265] = 16'h7c73;
    assign win_coe [266] = 16'h7c2b;
    assign win_coe [267] = 16'h7be1;
    assign win_coe [268] = 16'h7b93;
    assign win_coe [269] = 16'h7b44;
    assign win_coe [270] = 16'h7af1;
    assign win_coe [271] = 16'h7a9c;
    assign win_coe [272] = 16'h7a45;
    assign win_coe [273] = 16'h79ea;
    assign win_coe [274] = 16'h798e;
    assign win_coe [275] = 16'h792f;
    assign win_coe [276] = 16'h78cd;
    assign win_coe [277] = 16'h7869;
    assign win_coe [278] = 16'h7802;
    assign win_coe [279] = 16'h7799;
    assign win_coe [280] = 16'h772d;
    assign win_coe [281] = 16'h76bf;
    assign win_coe [282] = 16'h764e;
    assign win_coe [283] = 16'h75db;
    assign win_coe [284] = 16'h7566;
    assign win_coe [285] = 16'h74ef;
    assign win_coe [286] = 16'h7475;
    assign win_coe [287] = 16'h73f8;
    assign win_coe [288] = 16'h737a;
    assign win_coe [289] = 16'h72f9;
    assign win_coe [290] = 16'h7276;
    assign win_coe [291] = 16'h71f1;
    assign win_coe [292] = 16'h7169;
    assign win_coe [293] = 16'h70e0;
    assign win_coe [294] = 16'h7054;
    assign win_coe [295] = 16'h6fc6;
    assign win_coe [296] = 16'h6f36;
    assign win_coe [297] = 16'h6ea4;
    assign win_coe [298] = 16'h6e0f;
    assign win_coe [299] = 16'h6d79;
    assign win_coe [300] = 16'h6ce1;
    assign win_coe [301] = 16'h6c47;
    assign win_coe [302] = 16'h6bab;
    assign win_coe [303] = 16'h6b0d;
    assign win_coe [304] = 16'h6a6d;
    assign win_coe [305] = 16'h69cb;
    assign win_coe [306] = 16'h6927;
    assign win_coe [307] = 16'h6882;
    assign win_coe [308] = 16'h67da;
    assign win_coe [309] = 16'h6731;
    assign win_coe [310] = 16'h6687;
    assign win_coe [311] = 16'h65da;
    assign win_coe [312] = 16'h652c;
    assign win_coe [313] = 16'h647c;
    assign win_coe [314] = 16'h63cb;
    assign win_coe [315] = 16'h6318;
    assign win_coe [316] = 16'h6264;
    assign win_coe [317] = 16'h61ae;
    assign win_coe [318] = 16'h60f6;
    assign win_coe [319] = 16'h603d;
    assign win_coe [320] = 16'h5f83;
    assign win_coe [321] = 16'h5ec7;
    assign win_coe [322] = 16'h5e0a;
    assign win_coe [323] = 16'h5d4c;
    assign win_coe [324] = 16'h5c8c;
    assign win_coe [325] = 16'h5bcb;
    assign win_coe [326] = 16'h5b09;
    assign win_coe [327] = 16'h5a45;
    assign win_coe [328] = 16'h5981;
    assign win_coe [329] = 16'h58bb;
    assign win_coe [330] = 16'h57f4;
    assign win_coe [331] = 16'h572d;
    assign win_coe [332] = 16'h5664;
    assign win_coe [333] = 16'h559a;
    assign win_coe [334] = 16'h54cf;
    assign win_coe [335] = 16'h5404;
    assign win_coe [336] = 16'h5337;
    assign win_coe [337] = 16'h526a;
    assign win_coe [338] = 16'h519b;
    assign win_coe [339] = 16'h50cc;
    assign win_coe [340] = 16'h4ffd;
    assign win_coe [341] = 16'h4f2c;
    assign win_coe [342] = 16'h4e5b;
    assign win_coe [343] = 16'h4d89;
    assign win_coe [344] = 16'h4cb7;
    assign win_coe [345] = 16'h4be4;
    assign win_coe [346] = 16'h4b11;
    assign win_coe [347] = 16'h4a3d;
    assign win_coe [348] = 16'h4968;
    assign win_coe [349] = 16'h4894;
    assign win_coe [350] = 16'h47bf;
    assign win_coe [351] = 16'h46e9;
    assign win_coe [352] = 16'h4613;
    assign win_coe [353] = 16'h453d;
    assign win_coe [354] = 16'h4467;
    assign win_coe [355] = 16'h4390;
    assign win_coe [356] = 16'h42ba;
    assign win_coe [357] = 16'h41e3;
    assign win_coe [358] = 16'h410c;
    assign win_coe [359] = 16'h4035;
    assign win_coe [360] = 16'h3f5e;
    assign win_coe [361] = 16'h3e87;
    assign win_coe [362] = 16'h3db1;
    assign win_coe [363] = 16'h3cda;
    assign win_coe [364] = 16'h3c03;
    assign win_coe [365] = 16'h3b2d;
    assign win_coe [366] = 16'h3a57;
    assign win_coe [367] = 16'h3981;
    assign win_coe [368] = 16'h38ab;
    assign win_coe [369] = 16'h37d6;
    assign win_coe [370] = 16'h3701;
    assign win_coe [371] = 16'h362c;
    assign win_coe [372] = 16'h3558;
    assign win_coe [373] = 16'h3485;
    assign win_coe [374] = 16'h33b1;
    assign win_coe [375] = 16'h32df;
    assign win_coe [376] = 16'h320d;
    assign win_coe [377] = 16'h313b;
    assign win_coe [378] = 16'h306a;
    assign win_coe [379] = 16'h2f9a;
    assign win_coe [380] = 16'h2ecb;
    assign win_coe [381] = 16'h2dfc;
    assign win_coe [382] = 16'h2d2f;
    assign win_coe [383] = 16'h2c62;
    assign win_coe [384] = 16'h2b95;
    assign win_coe [385] = 16'h2aca;
    assign win_coe [386] = 16'h2a00;
    assign win_coe [387] = 16'h2937;
    assign win_coe [388] = 16'h286e;
    assign win_coe [389] = 16'h27a7;
    assign win_coe [390] = 16'h26e1;
    assign win_coe [391] = 16'h261c;
    assign win_coe [392] = 16'h2558;
    assign win_coe [393] = 16'h2495;
    assign win_coe [394] = 16'h23d3;
    assign win_coe [395] = 16'h2313;
    assign win_coe [396] = 16'h2254;
    assign win_coe [397] = 16'h2196;
    assign win_coe [398] = 16'h20da;
    assign win_coe [399] = 16'h201f;
    assign win_coe [400] = 16'h1f65;
    assign win_coe [401] = 16'h1ead;
    assign win_coe [402] = 16'h1df6;
    assign win_coe [403] = 16'h1d41;
    assign win_coe [404] = 16'h1c8d;
    assign win_coe [405] = 16'h1bdb;
    assign win_coe [406] = 16'h1b2b;
    assign win_coe [407] = 16'h1a7c;
    assign win_coe [408] = 16'h19ce;
    assign win_coe [409] = 16'h1923;
    assign win_coe [410] = 16'h1879;
    assign win_coe [411] = 16'h17d1;
    assign win_coe [412] = 16'h172a;
    assign win_coe [413] = 16'h1686;
    assign win_coe [414] = 16'h15e3;
    assign win_coe [415] = 16'h1542;
    assign win_coe [416] = 16'h14a3;
    assign win_coe [417] = 16'h1406;
    assign win_coe [418] = 16'h136b;
    assign win_coe [419] = 16'h12d2;
    assign win_coe [420] = 16'h123a;
    assign win_coe [421] = 16'h11a5;
    assign win_coe [422] = 16'h1112;
    assign win_coe [423] = 16'h1081;
    assign win_coe [424] = 16'h0ff2;
    assign win_coe [425] = 16'h0f65;
    assign win_coe [426] = 16'h0eda;
    assign win_coe [427] = 16'h0e52;
    assign win_coe [428] = 16'h0dcb;
    assign win_coe [429] = 16'h0d47;
    assign win_coe [430] = 16'h0cc5;
    assign win_coe [431] = 16'h0c46;
    assign win_coe [432] = 16'h0bc8;
    assign win_coe [433] = 16'h0b4d;
    assign win_coe [434] = 16'h0ad4;
    assign win_coe [435] = 16'h0a5e;
    assign win_coe [436] = 16'h09ea;
    assign win_coe [437] = 16'h0978;
    assign win_coe [438] = 16'h0909;
    assign win_coe [439] = 16'h089c;
    assign win_coe [440] = 16'h0832;
    assign win_coe [441] = 16'h07ca;
    assign win_coe [442] = 16'h0764;
    assign win_coe [443] = 16'h0701;
    assign win_coe [444] = 16'h06a1;
    assign win_coe [445] = 16'h0643;
    assign win_coe [446] = 16'h05e7;
    assign win_coe [447] = 16'h058e;
    assign win_coe [448] = 16'h0538;
    assign win_coe [449] = 16'h04e4;
    assign win_coe [450] = 16'h0493;
    assign win_coe [451] = 16'h0445;
    assign win_coe [452] = 16'h03f9;
    assign win_coe [453] = 16'h03b0;
    assign win_coe [454] = 16'h0369;
    assign win_coe [455] = 16'h0325;
    assign win_coe [456] = 16'h02e4;
    assign win_coe [457] = 16'h02a5;
    assign win_coe [458] = 16'h026a;
    assign win_coe [459] = 16'h0231;
    assign win_coe [460] = 16'h01fa;
    assign win_coe [461] = 16'h01c7;
    assign win_coe [462] = 16'h0196;
    assign win_coe [463] = 16'h0168;
    assign win_coe [464] = 16'h013c;
    assign win_coe [465] = 16'h0113;
    assign win_coe [466] = 16'h00ee;
    assign win_coe [467] = 16'h00cb;
    assign win_coe [468] = 16'h00aa;
    assign win_coe [469] = 16'h008d;
    assign win_coe [470] = 16'h0072;
    assign win_coe [471] = 16'h005a;
    assign win_coe [472] = 16'h0045;
    assign win_coe [473] = 16'h0033;
    assign win_coe [474] = 16'h0023;
    assign win_coe [475] = 16'h0017;
    assign win_coe [476] = 16'h000d;
    assign win_coe [477] = 16'h0006;
    assign win_coe [478] = 16'h0001;
    assign win_coe [479] = 16'h0000;

endmodule