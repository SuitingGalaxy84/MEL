`timescale 1ns / 1ps

module cpu_top #(
    parameter DATA_WIDTH = 32,
    parameter BOOT_ADDR = 32'h00000000
)(
    // ?��????????
    input  wire        clk,
    input  wire        rst_n,
    input  wire [31:0] if_id_instruction,
    
    // ?????????��?????��??��?????????????
    output wire [31:0] imem_addr,
    
    // === ?��???????????? ===
    output wire [31:0] debug_wb_data,    // WB?��????????
    output wire [4:0]  debug_wb_rd       // ?????????��??
);

// ================================================================
// ?????????��??
// ================================================================

// PC?��??????
wire [31:0] pc_out;
//wire [31:0] pc_plus_4;
wire [1:0]  pc_src; // ??��???????????PC????????


// ID?��??????????
wire [31:0] id_data1;
wire [31:0] id_data2;
wire [31:0] id_imm;

reg [31:0] id_ex_imm;

//reg        id_ex_alu_src_b;
//reg        id_ex_reg_write;

// EX/MEM?��?????????��?��??ALU?��????ALU?????????????��??????????????
reg [4:0]  ex_mem_rd;

wire [31:0] ex_mem_alu_result; // ??ALU??????????reg?��??

//reg        mem_wb_reg_write;
wire [4:0] ex_rd_out;

// ????????????????
wire        reg_write;
wire        alu_src_b;
wire        imm_control;
wire [3:0]  alu_control;
wire        forward_a;
wire        forward_b;

// ALU??����???��????��??��??????
wire        alu_zero_flag;

//adder 
wire [31:0] JumpTarget_Addr;

// ================================================================
// ???��??????
// ================================================================

// ???��?????��?��????????????????
Program_Counter pc_inst (
    .clk(clk),
    .reset_n(rst_n),
    .PC_Ctrl(pc_src),
    .JumpTarget_Addr(JumpTarget_Addr), // ��??��/??��???����
    .Boot_Addr(BOOT_ADDR),
    .PC_Out(pc_out)
//    .PC_Plus_4(pc_plus_4)
);

// ?????????????��???????��????
inst_decode #(
    .DATA_WIDTH(DATA_WIDTH)
) id_inst (
    .clk(clk),
    .rstn(rst_n),
    .sz_ext_select(imm_control),
    .we(reg_write),
    .data_in(ex_mem_alu_result), // ?????????��????��?ALU?��??
    .inst(if_id_instruction),
    .rd(ex_rd_out),
    .data1_pip(id_data1),
    .data2_pip(id_data2),
    .imm_gen_pip(id_imm)
);

// ?????????????��?��???��??????ex_mem_alu_result??
ALU #(
    .DW(DATA_WIDTH)
) alu_inst (
    .clk(clk),
    .rst_n(rst_n),
    .D1(id_data1),
    .D2(id_data2),
    .IG(id_ex_imm),
    .forward_a(forward_a),  // ???????��??
    .forward_b(forward_b),  // ???????��??
    .src_b(alu_src_b),
    .OP_ALU({2'b00, alu_control}), // ??????6??
    .R(ex_mem_alu_result), // ?��??????EX/MEM??ALU?��??
    .zero(alu_zero_flag)
);

//adder
Adder add_inst (
    .clk(clk),      // 50 MHz 
    .IG(id_ex_imm),
    .PCAD(pc_out),     
    .PCNAD(JumpTarget_Addr)     
);

// ????????
ControlUnit ctrl_inst (
    .clk(clk),
    .reset(!rst_n),
    .ins(if_id_instruction),
    .zero_flag(alu_zero_flag),
    .pc_src(pc_src) // ????PC????????
);

// delay
ControlSignalDelayer ctrlD_inst (
    .clk(clk),
    .reset(!rst_n),
    .reg_write_out(reg_write),
    .alu_src_b_out(alu_src_b),
    .imm_control_out(imm_control),
    .alu_control_out(alu_control),
    .ex_rd_out(ex_rd_out),
    .forward_a_out(forward_a),  // ?????��???����??��?????????��????
    .forward_b_out(forward_b)
);

// ================================================================
// ????
// ================================================================

// ???????��????
assign imem_addr = pc_out;

// WB?��??????
assign debug_wb_data = ex_mem_alu_result;
assign debug_wb_rd   = ex_rd_out;

endmodule